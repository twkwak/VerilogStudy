`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/03/24 18:49:33
// Design Name: 
// Module Name: tb_reg4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_reg4(
    input [3:0] data_in,
    input inen,
    input oen,
    input clk,
    input clr,
    input [3:0] data_out
    );
endmodule
