`timescale 1ns / 1ps
module control_block(z_f,s_f,clk,clr,opcode,pc_oen,mar_inen,rom_en,mdr_inen,     
    pc_inc,mdr_oen,ir_inen,tmp_inen,tmp_oen,creg_inen,creg_oen, 
    dreg_inen, dreg_oen,rreg_inen,rreg_oen,breg_inen,inreg_oen,keych_oen,
    outreg_inen, keyout_inen, load_pc,acc_oen,ah_inen,ah_reset,adds,subs,    
    ands,divs,muls,hs,ls);
    input [7:0] opcode; //명령어 입력
    input z_f,s_f,clk,clr;  //ALU의 계산 결과로 나오는 flag와 clk, clr
    output pc_oen,mar_inen,rom_en,mdr_inen,pc_inc,mdr_oen,ir_inen,tmp_inen,
             tmp_oen,creg_inen,creg_oen,dreg_inen,dreg_oen,rreg_inen, rreg_oen, 
             breg_inen,inreg_oen,keych_oen,outreg_inen,keyout_inen,
             load_pc,acc_oen,ah_inen,ah_reset,adds,subs,ands,divs,muls;
     output [1:0] hs,ls; //output의 전체 33개 신호는 각종 레지스터들의 최종 입출력 제어신호
     wire [11:0] t;        //ringcnt.v와 ctrl_signal.v 블록 연결을 위한 선
//decoder.v의 출력과 ctrl_signal.v 입력의 연결선
wire nop,outb,outs,add_s,sub_s,and_s, div_s,mul_s,shl,clr_s,psah,shr,load, jz,jmp,jge, mov_ah_cr, mov_ah_dr, mov_tmp_ah,mov_tmp_br,mov_tmp_cr, mov_tmp_dr,mov_tmp_rr,
     mov_cr_ah,mov_cr_br,mov_dr_ah, 
     mov_dr_tmp,mov_dr_br,mov_rr_ah,
     mov_key_ah,mov_inr_tmp,mov_inr_rr; 
  ringCounter u0(.clk(clk), .clr(clr), .t(t));  
  decoder u1(.ir_in(opcode),
            .nop(nop),
            .outb(outb),
            .outs(outs),
            .add_s(add_s),
            .sub_s(sub_s),
            .and_s(and_s),
            .div_s(div_s),
            .mul_s(mul_s),
            .shl(shl),
            .clr_s(clr_s),
            .psah(psah),
            .shr(shr),
            .load(load),
            .jz(jz),
            .jmp(jmp),
            .jge(jge),
            .mov_ah_cr(mov_ah_cr),
            .mov_ah_dr(mov_ah_dr),
            .mov_tmp_ah(mov_tmp_ah),
            .mov_tmp_br(mov_tmp_br),
            .mov_tmp_cr(mov_tmp_cr),
            .mov_tmp_dr(mov_tmp_dr),
            .mov_tmp_rr(mov_tmp_rr),
            .mov_cr_ah(mov_cr_ah),
            .mov_cr_br(mov_cr_br),
            .mov_dr_ah(mov_dr_ah),
            .mov_dr_tmp(mov_dr_tmp),
            .mov_dr_br(mov_dr_br),
            .mov_rr_ah(mov_rr_ah),
            .mov_key_ah(mov_key_ah),
            .mov_inr_tmp(mov_inr_tmp),
            .mov_inr_rr(mov_inr_rr)
            );

      control_signal u2(.t(t),
            .s_flag(s_f),
            .z_flag(z_f),
            .nop(nop),
            .outb(outb),
            .outs(outs),
            .add_s(add_s),
            .sub_s(sub_s),
            .and_s(and_s),
            .div_s(div_s),
            .mul_s(mul_s),
            .shl(shl),
            .clr_s(clr_s),
            .psah(psah),
            .shr(shr),
            .load(load),
            .jz(jz),
            .jmp(jmp),
            .jge(jge),
            .mov_ah_cr(mov_ah_cr),
            .mov_ah_dr(mov_ah_dr),
            .mov_tmp_ah(mov_tmp_ah),
            .mov_tmp_br(mov_tmp_br),
            .mov_tmp_cr(mov_tmp_cr),
            .mov_tmp_dr(mov_tmp_dr),
            .mov_tmp_rr(mov_tmp_rr),
            .mov_cr_ah(mov_cr_ah),
            .mov_cr_br(mov_cr_br),
            .mov_dr_ah(mov_dr_ah),
            .mov_dr_tmp(mov_dr_tmp),
            .mov_dr_br(mov_dr_br),
            .mov_rr_ah(mov_rr_ah),
            .mov_key_ah(mov_key_ah),
            .mov_inr_tmp(mov_inr_tmp),
            .mov_inr_rr(mov_inr_rr),
            .pc_oen(pc_oen),
            .mar_inen(mar_inen),
            .rom_en(rom_en),
            .mdr_inen(mdr_inen),
            .pc_inc(pc_inc),
            .mdr_oen(mdr_oen),
            .ir_inen(ir_inen),
            .tmp_inen(tmp_inen),
            .tmp_oen(tmp_oen),
            .creg_inen(creg_inen),
            .creg_oen(creg_oen),
            .dreg_inen(dreg_inen),
            .dreg_oen(dreg_oen),
            .rreg_inen(rreg_inen),
            .rreg_oen(rreg_oen),
            .breg_inen(breg_inen),
            .inreg_oen(inreg_oen),
            .keych_oen(keych_oen),
            .outreg_inen(outreg_inen),
            .keyout_inen(keyout_inen),
            .load_pc(load_pc),
            .acc_oen(acc_oen),
            .ah_inen(ah_inen),
            .ah_reset(ah_reset),
            .adds(adds),
            .subs(subs),
            .ands(ands),.divs(divs),
            .muls(muls), .hs(hs),
            .ls(ls)     );
  endmodule 
