`timescale 1ns/1ps

module tb_rv_fifo_1deep;

  localparam int DW = 32;

  // DUT I/O
  logic clk, rst_n;

  logic           in_valid;
  logic           in_ready;
  logic [DW-1:0]  in_data;

  logic           out_valid;
  logic           out_ready;
  logic [DW-1:0]  out_data;

  // Instantiate DUT
  rv_fifo_1deep #(.DW(DW)) dut (
    .clk(clk),
    .rst_n(rst_n),
    .in_valid(in_valid),
    .in_ready(in_ready),
    .in_data(in_data),
    .out_valid(out_valid),
    .out_ready(out_ready),
    .out_data(out_data)
  );

  // clock
  initial clk = 1'b0;
  always #5 clk = ~clk;

  // handshake events
  logic push, pop;
  assign push = in_valid  & in_ready;
  assign pop  = out_valid & out_ready;

  // reference model (1-depth)
  logic           ref_full;
  logic [DW-1:0]  ref_data;

  // stimulus control
  logic run_random;
  int unsigned next_payload;
  int unsigned cycle;

  // -----------------------
  // Reset task
  // -----------------------
  task automatic do_reset();
    begin
      rst_n = 1'b0;

      // TB-driven signals init
      in_valid    = 1'b0;       // one-bit zero
      in_data     = '0;         // all of bits are zero
      out_ready   = 1'b0;

      // REF init
      ref_full    = 1'b0;
      ref_data    = '0;

      // counters
      next_payload = 0;
      run_random   = 1'b0;

      repeat (3) @(posedge clk);
      rst_n = 1'b1;
      @(posedge clk);
    end
  endtask

  // -----------------------
  // Assertions (�ʼ� 2��)
  // -----------------------
  // stall ���� out_data ���� (���� ����Ŭ �������� üũ)
  assert property (@(posedge clk) disable iff (!rst_n)                  //assert ���ǿ� ���ÿ� ���� , �������̸� ���� x
    (out_valid && !out_ready) |=> (out_data == $past(out_data))     //need to hold data when out_valid= 1 && out_ready = 0 , |=> ����Ŭ������ ��ȭ
  ) else $fatal(1, "out_data changed while stalled");


  // out_valid�� accept(pop)�� ������ ����
  assert property (@(posedge clk) disable iff (!rst_n)
    (out_valid && !out_ready) |=> out_valid                         //out_valid must be 1 at next cycle
  ) else $fatal(1, "out_valid dropped before acceptance");

  // -----------------------
  // ������ ����̹�: negedge������ stimulus ����
  // (��Ƽ����̺� ����)
  // -----------------------
  always @(negedge clk) begin
    if (!rst_n) begin
      out_ready <= 1'b0;
      in_valid  <= 1'b0;
      in_data   <= '0;
    end 
    else if (run_random)                    //random value ���� �� push �߻� �� data update
    begin
      // random backpressure
      out_ready <= $urandom_range(0,1);

      // random valid (70% Ȯ��)
      in_valid  <= ($urandom_range(0,99) < 70);

      // sender rule: push�� ���� data ����
    if (in_valid && in_ready) 
      begin       //push!
        in_data <= next_payload[DW-1:0];    //   data update at negedge && push
      end
      // else: in_data ���� (stall ���� data stable)
    end 
    
    else // 300 cycle end , run_random = 0 
    begin
      // drain mode
      out_ready <= 1'b1;
      in_valid  <= 1'b0;
      // in_data�� �ǹ� ����(��ȿ �ƴ�) -> �״�� �ֵ� ��
    end
  end

  // -----------------------
  // Reference model + checking (posedge����)
  // -----------------------
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      ref_full <= 1'b0;
      ref_data <= '0;
    end else begin
      // pop �߻� �� ������ üũ pop = out_valid= 1 , out_ready= 1, full= 1�϶� �߻�
      if (pop) 
      begin
        if (!ref_full) $fatal(1, "REF underflow: pop but ref_full=0");              // pop���� full=0 �� ����
        if (out_data !== ref_data) $fatal(1, "DATA mismatch: exp=0x%08h got=0x%08h", ref_data, out_data);       
      end

      // ref ���� ������Ʈ
      unique case ({push, pop})
        2'b10: begin // push only
          if (ref_full) $fatal(1, "REF overflow: push but ref_full=1");
          ref_data <= in_data;
          ref_full <= 1'b1;
          next_payload <= next_payload + 1;
        end
        2'b01: begin // pop only
          ref_full <= 1'b0;
        end
        2'b11: begin // push & pop
          ref_data <= in_data;  // replace with new
          ref_full <= 1'b1;
          next_payload <= next_payload + 1;
        end
        default: ; // no event
      endcase
    end
  end

  // -----------------------
  // Main test sequence
  // -----------------------
  initial begin
    do_reset();

    // 1) random test phase
    run_random = 1'b1;
    for (cycle = 0; cycle < 300; cycle++) begin
      @(posedge clk);
    end

    // 2) drain phase
    run_random = 1'b0;
    repeat (20) @(posedge clk);

    // drain Ȯ��: DUT�� REF �� �� ���� ��
    if (out_valid) $fatal(1, "Drain failed: DUT still valid");
    if (ref_full)  $fatal(1, "Drain failed: ref_full still 1");

    $display("PASS ? Project 1 TB complete");
    $finish;
  end

endmodule